* C:\Projekte\20171122 Maxima Thermal Modeling\coupled-thermal-resistor-model.asc
R1 n5 n1 0.05
R2 n2 n6 0.1
R3 n7 n3 0.075
R4 n8 n4 0.1
R5 0 n5 0.1
R6 n6 0 0.1
R7 n7 0 0.1
R8 0 n8 0.1
R9 n5 n6 1
R10 n7 n6 0.5
R11 n7 n8 1
R12 n8 n5 0.5
R13 n5 n7 2
R14 n8 n6 2
I1 0 n1 1
I2 0 n2 0
I3 0 n3 0
I4 0 n4 0
I5 n2 n4 0
V1 n6 n8 0
C1 n5 n8 1
L1 n0 n4 1
.end


